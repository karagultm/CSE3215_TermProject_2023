module cpu ();




endmodule