module d_latch (
    input D, C;
    output Q;
    wire R, S1 , R1 ;


);
    
endmodule